module CPU();

reg [63:0] IR, [63:0] PC;
reg [63:0] MAR, [63:0] MDR;




endmodule