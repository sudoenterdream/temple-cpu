module ControlUnit();


endmodule